
module gaming
	(
		CLOCK_50,						//	On Board 50 MHz
		// Your inputs and outputs here
		KEY,		
		SW,// On Board Keys
		// The ports below are for the VGA output.  Do not change.
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B   						//	VGA Blue[9:0]
	);

	input			CLOCK_50;				//	50 MHz
	input	[3:0]	KEY;		
	input [9:0] SW;
	// Declare your inputs and outputs here
	// Do not change the following outputs
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK_N;				//	VGA BLANK
	output			VGA_SYNC_N;				//	VGA SYNC
	output	[7:0]	VGA_R;   				//	VGA Red[7:0] Changed from 10 to 8-bit DAC
	output	[7:0]	VGA_G;	 				//	VGA Green[7:0]
	output	[7:0]	VGA_B;   				//	VGA Blue[7:0]
	
	wire resetn;
	assign resetn = KEY[0];
	
	// Create the colour, x, y and writeEn wires that are inputs to the controller.

	wire [2:0] colour;
	wire [8:0] x;
	wire [7:0] y;
	wire writeEn;

	// Create an Instance of a VGA controller - there can be only one!
	// Define the number of colours as well as the initial background
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(colour),
			.x(x),
			.y(y),
			.plot(1'b1),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK_N),
			.VGA_SYNC(VGA_SYNC_N),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "320x240";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "black.mif";
			
	wire L_x, L_y, L_c,plot_enable, black_enable, done;
	assign resetn = KEY[0];
				
	Counter U2(resetn, CLOCK_50,x,y);
	vga_pic U1(CLOCK_50, resetn, x,y,colour);
					
endmodule


module vga_pic(
input wire clk , 
input wire reset , 
input wire [8:0] x , //x coordinate
input wire [7:0] y , //y coordinate

output reg [2:0] colour//output color
);

parameter x_initial= 10'd122,  //begins at  
y_initial= 10'd0 ; //begins at

parameter width = 10'd76,  //width  should be able be divided by four 
height = 10'd240 ; //height


wire [6:0] char_x ; //x coordinate 0-89
wire [7:0] char_y ; //y coordinate 0-239


//Check if it reaches the area of title
assign char_x = (((x >= x_initial) && (x < (x_initial + width)))
&&((y >= y_initial)&&(y < (y_initial + height))))
? (x - x_initial) : 0;

assign char_y = (((x >= x_initial) && (x < (x_initial + width)))
&&((y >= y_initial)&&(y < (y_initial + height))))
? (y - y_initial) : 0;

//reg [89:0] initial_value = 90'h80000300000C0000300001;
//char:Title 
reg [75:0] char [239:0]; //Title LCD character font
always@(*)
begin
	 char[0]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[1]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[2]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[3]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[4]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[5]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[6]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[7]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[8]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[9]  <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[10] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[11] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[12] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[13] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[14] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[15] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[16] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[17] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[18] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[19] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[20] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[21] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[22] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[23] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[24] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[25] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[26] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[27] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[28] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[29] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[30] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[31] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[32] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[33] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[34] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[35] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[36] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[37] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[38] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[39] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[40] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[41] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[42] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[43] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[44] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[45] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[46] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[47] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[48] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[49] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[50] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[51] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[52] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[53] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[54] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[55] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[56] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[57] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[58] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[59] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[60] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[61] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[62] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[63] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[64] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[65] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[66] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[67] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[68] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[69] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[70] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[71] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[72] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[73] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[74] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[75] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[76] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[77] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[78] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[79] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[80] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[81] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[82] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[83] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[84] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[85] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[86] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[87] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[88] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[89] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[90] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[91] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[92] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[93] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[94] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[95] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[96] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[97] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[98] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[99] <= 76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[100] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[101] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[102] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[103] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[104] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[105] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[106] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[107] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[108] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[109] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[110] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[111] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[112] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[113] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[114] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[115] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[116] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[117] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[118] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[119] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[120] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[121] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[122] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[123] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[124] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[125] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[126] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[127] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[128] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[129] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[130] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[131] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[132] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[133] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[134] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[135] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[136] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[137] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[138] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[139] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[140] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[141] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[142] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[143] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[144] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[145] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[146] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[147] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[148] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[149] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[150] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[151] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[152] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[153] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[154] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[155] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[156] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[157] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[158] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[159] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[160] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[161] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[162] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[163] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[164] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[165] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[166] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[167] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[168] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[169] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[170] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[171] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[172] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[173] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[174] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[175] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[176] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[177] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[178] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[179] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[180] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[181] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[182] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[183] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[184] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[185] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[186] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[187] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[188] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[189] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[190] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[191] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[192] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[193] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[194] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[195] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[196] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[197] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[198] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[199] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[200] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[201] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[202] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[203] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[204] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[205] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[206] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[207] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[208] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[209] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[210] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[211] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[212] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[213] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[214] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[215] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[216] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[217] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[218] <=76'b0011111111111111111111111111111111111111111111111111111111111111111111111111;
    char[219] <=76'b0011111111111111111111111111111111111111111111111111111111111111111111111111;
    char[220] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[221] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[222] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[223] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[224] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[225] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[226] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[227] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[228] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[229] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[230] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[231] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[232] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[233] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[234] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[235] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[236] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[237] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[238] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
    char[239] <=76'b0011000000000000000011000000000000000011000000000000000011000000000000000011;
end

 always@(posedge clk or negedge reset)
 if(!reset)
 colour <= 3'b111;
 
 else if((((x >= (x_initial - 1'b1))
 && (x < (x_initial + width -1'b1)))
 && ((y >= y_initial) && (y < (y_initial + height))))
 && (char[char_y][10'd74 - char_x] == 1'b1))
 colour <= 3'b000;
 else
 colour <= 3'b111;

endmodule


module Counter(reset,clk,xout, yout);
input reset,clk;
output reg [8:0] xout;
output reg[7:0] yout;
reg [16:0] counter;

always@(posedge clk)
begin
	if(!reset)
	begin
		counter <=0;
	end
	else 
	begin
		if (counter == 17'b11111111111111111)
		begin
			xout <= counter[8:0];
			yout <= counter[16:9];
			counter <= 17'b0;
		end
		else
		begin
		counter <= counter + 1;
		xout <= counter[8:0];
		yout <= counter[16 :9];
		end
	end
end

endmodule
